`include "uart.sv"
`include "uart_rx.sv"
`include "uart_tx.sv"

`include "tb_uart_top.sv"

